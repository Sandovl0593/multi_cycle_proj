module extend (
    input wire [23:0] Instr,
    input wire [1:0] ImmSrc,
    output reg [31:0] ExtImm
);
    always @(*)
        case (ImmSrc)
            2'b00: ExtImm =  ({24'b000000000000000000000000, Instr[7:0]}>>2*Instr[11:8]) |
                             ({24'b000000000000000000000000, Instr[7:0]}<<32-2*Instr[11:8]); // Zero-extend para DP with rota
            2'b01: ExtImm = {20'b00000000000000000000, Instr[11:0]};     // Zero-extend para Load/Store
            2'b10: ExtImm = {{6 {Instr[23]}}, Instr[23:0], 2'b00};       // Sign-extend para Branch
            default: ExtImm = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
        endcase
endmodule